// =============================================================================
// Filename: glitch_free.v
// Author: KANG, Jian
// Email: jkangac@connect.ust.hk
// Affiliation: Hong Kong University of Science and Technology
// Description:
// -----------------------------------------------------------------------------
`timescale 1 ns / 1 ps
module glitch_free(
	input clk,
	input rst,
		
);

endmodule